module LDST_KFMMC_SPI2IDE_ROM (clock, address, data_out);
    input clock;
    input [10:0] address;
    output reg [12:0] data_out;

    always @ (posedge clock)
    begin
        case (address)
            11'h0000: data_out = 12'h203;
            11'h0001: data_out = 12'h182;
            11'h0002: data_out = 12'h280;
            11'h0003: data_out = 12'h1c3;
            11'h0004: data_out = 12'h200;
            11'h0005: data_out = 12'h1c4;
            11'h0006: data_out = 12'h20a;
            11'h0007: data_out = 12'h104;
            11'h0008: data_out = 12'h2ff;
            11'h0009: data_out = 12'h180;
            11'h000a: data_out = 12'h205;
            11'h000b: data_out = 12'h4f0;
            11'h000c: data_out = 12'h004;
            11'h000d: data_out = 12'h100;
            11'h000e: data_out = 12'h201;
            11'h000f: data_out = 12'h101;
            11'h0010: data_out = 12'h282;
            11'h0011: data_out = 12'h103;
            11'h0012: data_out = 12'h003;
            11'h0013: data_out = 12'h104;
            11'h0014: data_out = 12'h200;
            11'h0015: data_out = 12'h918;
            11'h0016: data_out = 12'h200;
            11'h0017: data_out = 12'h808;
            11'h0018: data_out = 12'h2fd;
            11'h0019: data_out = 12'h100;
            11'h001a: data_out = 12'h205;
            11'h001b: data_out = 12'h4db;
            11'h001c: data_out = 12'h240;
            11'h001d: data_out = 12'h180;
            11'h001e: data_out = 12'h205;
            11'h001f: data_out = 12'h4f0;
            11'h0020: data_out = 12'h206;
            11'h0021: data_out = 12'h40d;
            11'h0022: data_out = 12'h295;
            11'h0023: data_out = 12'h180;
            11'h0024: data_out = 12'h205;
            11'h0025: data_out = 12'h4f0;
            11'h0026: data_out = 12'h20a;
            11'h0027: data_out = 12'h104;
            11'h0028: data_out = 12'h206;
            11'h0029: data_out = 12'h41e;
            11'h002a: data_out = 12'h005;
            11'h002b: data_out = 12'h100;
            11'h002c: data_out = 12'h201;
            11'h002d: data_out = 12'h101;
            11'h002e: data_out = 12'h240;
            11'h002f: data_out = 12'h103;
            11'h0030: data_out = 12'h003;
            11'h0031: data_out = 12'h200;
            11'h0032: data_out = 12'h935;
            11'h0033: data_out = 12'h200;
            11'h0034: data_out = 12'h800;
            11'h0035: data_out = 12'h082;
            11'h0036: data_out = 12'h100;
            11'h0037: data_out = 12'h204;
            11'h0038: data_out = 12'h101;
            11'h0039: data_out = 12'h200;
            11'h003a: data_out = 12'h103;
            11'h003b: data_out = 12'h003;
            11'h003c: data_out = 12'h200;
            11'h003d: data_out = 12'h963;
            11'h003e: data_out = 12'h2ff;
            11'h003f: data_out = 12'h106;
            11'h0040: data_out = 12'h241;
            11'h0041: data_out = 12'h180;
            11'h0042: data_out = 12'h205;
            11'h0043: data_out = 12'h4f0;
            11'h0044: data_out = 12'h205;
            11'h0045: data_out = 12'h4fc;
            11'h0046: data_out = 12'h2f9;
            11'h0047: data_out = 12'h180;
            11'h0048: data_out = 12'h205;
            11'h0049: data_out = 12'h4f0;
            11'h004a: data_out = 12'h20a;
            11'h004b: data_out = 12'h104;
            11'h004c: data_out = 12'h206;
            11'h004d: data_out = 12'h41e;
            11'h004e: data_out = 12'h005;
            11'h004f: data_out = 12'h100;
            11'h0050: data_out = 12'h200;
            11'h0051: data_out = 12'h101;
            11'h0052: data_out = 12'h240;
            11'h0053: data_out = 12'h103;
            11'h0054: data_out = 12'h003;
            11'h0055: data_out = 12'h200;
            11'h0056: data_out = 12'h9e6;
            11'h0057: data_out = 12'h006;
            11'h0058: data_out = 12'h100;
            11'h0059: data_out = 12'h201;
            11'h005a: data_out = 12'h101;
            11'h005b: data_out = 12'h282;
            11'h005c: data_out = 12'h103;
            11'h005d: data_out = 12'h003;
            11'h005e: data_out = 12'h106;
            11'h005f: data_out = 12'h200;
            11'h0060: data_out = 12'h900;
            11'h0061: data_out = 12'h200;
            11'h0062: data_out = 12'h840;
            11'h0063: data_out = 12'h206;
            11'h0064: data_out = 12'h408;
            11'h0065: data_out = 12'h248;
            11'h0066: data_out = 12'h180;
            11'h0067: data_out = 12'h205;
            11'h0068: data_out = 12'h4f0;
            11'h0069: data_out = 12'h200;
            11'h006a: data_out = 12'h180;
            11'h006b: data_out = 12'h205;
            11'h006c: data_out = 12'h4f0;
            11'h006d: data_out = 12'h200;
            11'h006e: data_out = 12'h180;
            11'h006f: data_out = 12'h205;
            11'h0070: data_out = 12'h4f0;
            11'h0071: data_out = 12'h201;
            11'h0072: data_out = 12'h180;
            11'h0073: data_out = 12'h205;
            11'h0074: data_out = 12'h4f0;
            11'h0075: data_out = 12'h2aa;
            11'h0076: data_out = 12'h180;
            11'h0077: data_out = 12'h205;
            11'h0078: data_out = 12'h4f0;
            11'h0079: data_out = 12'h287;
            11'h007a: data_out = 12'h180;
            11'h007b: data_out = 12'h205;
            11'h007c: data_out = 12'h4f0;
            11'h007d: data_out = 12'h20a;
            11'h007e: data_out = 12'h104;
            11'h007f: data_out = 12'h206;
            11'h0080: data_out = 12'h41e;
            11'h0081: data_out = 12'h005;
            11'h0082: data_out = 12'h100;
            11'h0083: data_out = 12'h201;
            11'h0084: data_out = 12'h101;
            11'h0085: data_out = 12'h240;
            11'h0086: data_out = 12'h103;
            11'h0087: data_out = 12'h003;
            11'h0088: data_out = 12'h200;
            11'h0089: data_out = 12'h990;
            11'h008a: data_out = 12'h204;
            11'h008b: data_out = 12'h100;
            11'h008c: data_out = 12'h205;
            11'h008d: data_out = 12'h4d4;
            11'h008e: data_out = 12'h200;
            11'h008f: data_out = 12'h806;
            11'h0090: data_out = 12'h206;
            11'h0091: data_out = 12'h400;
            11'h0092: data_out = 12'h080;
            11'h0093: data_out = 12'h100;
            11'h0094: data_out = 12'h201;
            11'h0095: data_out = 12'h101;
            11'h0096: data_out = 12'h200;
            11'h0097: data_out = 12'h103;
            11'h0098: data_out = 12'h003;
            11'h0099: data_out = 12'h200;
            11'h009a: data_out = 12'h900;
            11'h009b: data_out = 12'h2ff;
            11'h009c: data_out = 12'h180;
            11'h009d: data_out = 12'h205;
            11'h009e: data_out = 12'h4f0;
            11'h009f: data_out = 12'h080;
            11'h00a0: data_out = 12'h100;
            11'h00a1: data_out = 12'h2aa;
            11'h00a2: data_out = 12'h101;
            11'h00a3: data_out = 12'h282;
            11'h00a4: data_out = 12'h103;
            11'h00a5: data_out = 12'h003;
            11'h00a6: data_out = 12'h200;
            11'h00a7: data_out = 12'h9aa;
            11'h00a8: data_out = 12'h200;
            11'h00a9: data_out = 12'h800;
            11'h00aa: data_out = 12'h206;
            11'h00ab: data_out = 12'h408;
            11'h00ac: data_out = 12'h277;
            11'h00ad: data_out = 12'h180;
            11'h00ae: data_out = 12'h205;
            11'h00af: data_out = 12'h4f0;
            11'h00b0: data_out = 12'h206;
            11'h00b1: data_out = 12'h40d;
            11'h00b2: data_out = 12'h20a;
            11'h00b3: data_out = 12'h104;
            11'h00b4: data_out = 12'h206;
            11'h00b5: data_out = 12'h41e;
            11'h00b6: data_out = 12'h005;
            11'h00b7: data_out = 12'h100;
            11'h00b8: data_out = 12'h201;
            11'h00b9: data_out = 12'h101;
            11'h00ba: data_out = 12'h240;
            11'h00bb: data_out = 12'h103;
            11'h00bc: data_out = 12'h003;
            11'h00bd: data_out = 12'h200;
            11'h00be: data_out = 12'h9c1;
            11'h00bf: data_out = 12'h200;
            11'h00c0: data_out = 12'h800;
            11'h00c1: data_out = 12'h206;
            11'h00c2: data_out = 12'h408;
            11'h00c3: data_out = 12'h269;
            11'h00c4: data_out = 12'h180;
            11'h00c5: data_out = 12'h205;
            11'h00c6: data_out = 12'h4f0;
            11'h00c7: data_out = 12'h240;
            11'h00c8: data_out = 12'h180;
            11'h00c9: data_out = 12'h205;
            11'h00ca: data_out = 12'h4f0;
            11'h00cb: data_out = 12'h2ff;
            11'h00cc: data_out = 12'h180;
            11'h00cd: data_out = 12'h205;
            11'h00ce: data_out = 12'h4f0;
            11'h00cf: data_out = 12'h280;
            11'h00d0: data_out = 12'h180;
            11'h00d1: data_out = 12'h205;
            11'h00d2: data_out = 12'h4f0;
            11'h00d3: data_out = 12'h200;
            11'h00d4: data_out = 12'h180;
            11'h00d5: data_out = 12'h205;
            11'h00d6: data_out = 12'h4f0;
            11'h00d7: data_out = 12'h20a;
            11'h00d8: data_out = 12'h104;
            11'h00d9: data_out = 12'h206;
            11'h00da: data_out = 12'h41e;
            11'h00db: data_out = 12'h005;
            11'h00dc: data_out = 12'h100;
            11'h00dd: data_out = 12'h200;
            11'h00de: data_out = 12'h101;
            11'h00df: data_out = 12'h240;
            11'h00e0: data_out = 12'h103;
            11'h00e1: data_out = 12'h003;
            11'h00e2: data_out = 12'h200;
            11'h00e3: data_out = 12'h9e6;
            11'h00e4: data_out = 12'h200;
            11'h00e5: data_out = 12'h8aa;
            11'h00e6: data_out = 12'h206;
            11'h00e7: data_out = 12'h408;
            11'h00e8: data_out = 12'h249;
            11'h00e9: data_out = 12'h180;
            11'h00ea: data_out = 12'h205;
            11'h00eb: data_out = 12'h4f0;
            11'h00ec: data_out = 12'h206;
            11'h00ed: data_out = 12'h40d;
            11'h00ee: data_out = 12'h20a;
            11'h00ef: data_out = 12'h104;
            11'h00f0: data_out = 12'h206;
            11'h00f1: data_out = 12'h41e;
            11'h00f2: data_out = 12'h005;
            11'h00f3: data_out = 12'h100;
            11'h00f4: data_out = 12'h200;
            11'h00f5: data_out = 12'h101;
            11'h00f6: data_out = 12'h240;
            11'h00f7: data_out = 12'h103;
            11'h00f8: data_out = 12'h003;
            11'h00f9: data_out = 12'h200;
            11'h00fa: data_out = 12'h9fd;
            11'h00fb: data_out = 12'h200;
            11'h00fc: data_out = 12'h800;
            11'h00fd: data_out = 12'h20a;
            11'h00fe: data_out = 12'h104;
            11'h00ff: data_out = 12'h2fe;
            11'h0100: data_out = 12'h105;
            11'h0101: data_out = 12'h206;
            11'h0102: data_out = 12'h439;
            11'h0103: data_out = 12'h006;
            11'h0104: data_out = 12'h100;
            11'h0105: data_out = 12'h2fe;
            11'h0106: data_out = 12'h101;
            11'h0107: data_out = 12'h240;
            11'h0108: data_out = 12'h103;
            11'h0109: data_out = 12'h003;
            11'h010a: data_out = 12'h201;
            11'h010b: data_out = 12'h90e;
            11'h010c: data_out = 12'h200;
            11'h010d: data_out = 12'h800;
            11'h010e: data_out = 12'h210;
            11'h010f: data_out = 12'h104;
            11'h0110: data_out = 12'h2ff;
            11'h0111: data_out = 12'h180;
            11'h0112: data_out = 12'h205;
            11'h0113: data_out = 12'h4f0;
            11'h0114: data_out = 12'h080;
            11'h0115: data_out = 12'h185;
            11'h0116: data_out = 12'h004;
            11'h0117: data_out = 12'h100;
            11'h0118: data_out = 12'h201;
            11'h0119: data_out = 12'h101;
            11'h011a: data_out = 12'h282;
            11'h011b: data_out = 12'h103;
            11'h011c: data_out = 12'h003;
            11'h011d: data_out = 12'h104;
            11'h011e: data_out = 12'h201;
            11'h011f: data_out = 12'h922;
            11'h0120: data_out = 12'h201;
            11'h0121: data_out = 12'h810;
            11'h0122: data_out = 12'h206;
            11'h0123: data_out = 12'h408;
            11'h0124: data_out = 12'h27a;
            11'h0125: data_out = 12'h180;
            11'h0126: data_out = 12'h205;
            11'h0127: data_out = 12'h4f0;
            11'h0128: data_out = 12'h206;
            11'h0129: data_out = 12'h40d;
            11'h012a: data_out = 12'h20a;
            11'h012b: data_out = 12'h104;
            11'h012c: data_out = 12'h206;
            11'h012d: data_out = 12'h41e;
            11'h012e: data_out = 12'h005;
            11'h012f: data_out = 12'h100;
            11'h0130: data_out = 12'h200;
            11'h0131: data_out = 12'h101;
            11'h0132: data_out = 12'h240;
            11'h0133: data_out = 12'h103;
            11'h0134: data_out = 12'h003;
            11'h0135: data_out = 12'h201;
            11'h0136: data_out = 12'h939;
            11'h0137: data_out = 12'h200;
            11'h0138: data_out = 12'h800;
            11'h0139: data_out = 12'h2bf;
            11'h013a: data_out = 12'h100;
            11'h013b: data_out = 12'h205;
            11'h013c: data_out = 12'h4db;
            11'h013d: data_out = 12'h2ff;
            11'h013e: data_out = 12'h180;
            11'h013f: data_out = 12'h205;
            11'h0140: data_out = 12'h4f0;
            11'h0141: data_out = 12'h080;
            11'h0142: data_out = 12'h100;
            11'h0143: data_out = 12'h240;
            11'h0144: data_out = 12'h101;
            11'h0145: data_out = 12'h200;
            11'h0146: data_out = 12'h103;
            11'h0147: data_out = 12'h003;
            11'h0148: data_out = 12'h100;
            11'h0149: data_out = 12'h205;
            11'h014a: data_out = 12'h4d4;
            11'h014b: data_out = 12'h206;
            11'h014c: data_out = 12'h400;
            11'h014d: data_out = 12'h08c;
            11'h014e: data_out = 12'h104;
            11'h014f: data_out = 12'h08d;
            11'h0150: data_out = 12'h105;
            11'h0151: data_out = 12'h08e;
            11'h0152: data_out = 12'h106;
            11'h0153: data_out = 12'h08f;
            11'h0154: data_out = 12'h107;
            11'h0155: data_out = 12'h200;
            11'h0156: data_out = 12'h190;
            11'h0157: data_out = 12'h191;
            11'h0158: data_out = 12'h20f;
            11'h0159: data_out = 12'h192;
            11'h015a: data_out = 12'h23f;
            11'h015b: data_out = 12'h193;
            11'h015c: data_out = 12'h004;
            11'h015d: data_out = 12'h100;
            11'h015e: data_out = 12'h2b1;
            11'h015f: data_out = 12'h101;
            11'h0160: data_out = 12'h282;
            11'h0161: data_out = 12'h103;
            11'h0162: data_out = 12'h003;
            11'h0163: data_out = 12'h104;
            11'h0164: data_out = 12'h005;
            11'h0165: data_out = 12'h100;
            11'h0166: data_out = 12'h203;
            11'h0167: data_out = 12'h101;
            11'h0168: data_out = 12'h283;
            11'h0169: data_out = 12'h103;
            11'h016a: data_out = 12'h003;
            11'h016b: data_out = 12'h105;
            11'h016c: data_out = 12'h200;
            11'h016d: data_out = 12'h101;
            11'h016e: data_out = 12'h006;
            11'h016f: data_out = 12'h100;
            11'h0170: data_out = 12'h003;
            11'h0171: data_out = 12'h106;
            11'h0172: data_out = 12'h007;
            11'h0173: data_out = 12'h100;
            11'h0174: data_out = 12'h003;
            11'h0175: data_out = 12'h107;
            11'h0176: data_out = 12'h201;
            11'h0177: data_out = 12'ha7a;
            11'h0178: data_out = 12'h201;
            11'h0179: data_out = 12'h896;
            11'h017a: data_out = 12'h090;
            11'h017b: data_out = 12'h100;
            11'h017c: data_out = 12'h201;
            11'h017d: data_out = 12'h101;
            11'h017e: data_out = 12'h280;
            11'h017f: data_out = 12'h103;
            11'h0180: data_out = 12'h003;
            11'h0181: data_out = 12'h190;
            11'h0182: data_out = 12'h091;
            11'h0183: data_out = 12'h100;
            11'h0184: data_out = 12'h200;
            11'h0185: data_out = 12'h101;
            11'h0186: data_out = 12'h281;
            11'h0187: data_out = 12'h103;
            11'h0188: data_out = 12'h003;
            11'h0189: data_out = 12'h191;
            11'h018a: data_out = 12'h101;
            11'h018b: data_out = 12'h240;
            11'h018c: data_out = 12'h100;
            11'h018d: data_out = 12'h282;
            11'h018e: data_out = 12'h103;
            11'h018f: data_out = 12'h003;
            11'h0190: data_out = 12'h201;
            11'h0191: data_out = 12'ha5c;
            11'h0192: data_out = 12'h2ff;
            11'h0193: data_out = 12'h190;
            11'h0194: data_out = 12'h23f;
            11'h0195: data_out = 12'h191;
            11'h0196: data_out = 12'h090;
            11'h0197: data_out = 12'h194;
            11'h0198: data_out = 12'h091;
            11'h0199: data_out = 12'h195;
            11'h019a: data_out = 12'h092;
            11'h019b: data_out = 12'h196;
            11'h019c: data_out = 12'h093;
            11'h019d: data_out = 12'h197;
            11'h019e: data_out = 12'h2fe;
            11'h019f: data_out = 12'h100;
            11'h01a0: data_out = 12'h205;
            11'h01a1: data_out = 12'h4e9;
            11'h01a2: data_out = 12'h200;
            11'h01a3: data_out = 12'h1c4;
            11'h01a4: data_out = 12'h201;
            11'h01a5: data_out = 12'h1c6;
            11'h01a6: data_out = 12'h201;
            11'h01a7: data_out = 12'h1c7;
            11'h01a8: data_out = 12'h200;
            11'h01a9: data_out = 12'h1c8;
            11'h01aa: data_out = 12'h1c9;
            11'h01ab: data_out = 12'h1ca;
            11'h01ac: data_out = 12'h1cb;
            11'h01ad: data_out = 12'h204;
            11'h01ae: data_out = 12'h4fd;
            11'h01af: data_out = 12'h2fe;
            11'h01b0: data_out = 12'h100;
            11'h01b1: data_out = 12'h205;
            11'h01b2: data_out = 12'h4db;
            11'h01b3: data_out = 12'h27f;
            11'h01b4: data_out = 12'h100;
            11'h01b5: data_out = 12'h205;
            11'h01b6: data_out = 12'h4e9;
            11'h01b7: data_out = 12'h240;
            11'h01b8: data_out = 12'h100;
            11'h01b9: data_out = 12'h205;
            11'h01ba: data_out = 12'h4e2;
            11'h01bb: data_out = 12'h202;
            11'h01bc: data_out = 12'h181;
            11'h01bd: data_out = 12'h0c3;
            11'h01be: data_out = 12'h100;
            11'h01bf: data_out = 12'h280;
            11'h01c0: data_out = 12'h101;
            11'h01c1: data_out = 12'h200;
            11'h01c2: data_out = 12'h103;
            11'h01c3: data_out = 12'h003;
            11'h01c4: data_out = 12'h201;
            11'h01c5: data_out = 12'h9bd;
            11'h01c6: data_out = 12'h0cd;
            11'h01c7: data_out = 12'h100;
            11'h01c8: data_out = 12'h290;
            11'h01c9: data_out = 12'h101;
            11'h01ca: data_out = 12'h240;
            11'h01cb: data_out = 12'h103;
            11'h01cc: data_out = 12'h003;
            11'h01cd: data_out = 12'h201;
            11'h01ce: data_out = 12'h99e;
            11'h01cf: data_out = 12'h0cb;
            11'h01d0: data_out = 12'h100;
            11'h01d1: data_out = 12'h201;
            11'h01d2: data_out = 12'h101;
            11'h01d3: data_out = 12'h200;
            11'h01d4: data_out = 12'h103;
            11'h01d5: data_out = 12'h003;
            11'h01d6: data_out = 12'h201;
            11'h01d7: data_out = 12'h9af;
            11'h01d8: data_out = 12'h200;
            11'h01d9: data_out = 12'h1c4;
            11'h01da: data_out = 12'h2b6;
            11'h01db: data_out = 12'h100;
            11'h01dc: data_out = 12'h205;
            11'h01dd: data_out = 12'h4e9;
            11'h01de: data_out = 12'h240;
            11'h01df: data_out = 12'h103;
            11'h01e0: data_out = 12'h0cd;
            11'h01e1: data_out = 12'h100;
            11'h01e2: data_out = 12'h208;
            11'h01e3: data_out = 12'h101;
            11'h01e4: data_out = 12'h003;
            11'h01e5: data_out = 12'h200;
            11'h01e6: data_out = 12'h900;
            11'h01e7: data_out = 12'h291;
            11'h01e8: data_out = 12'h101;
            11'h01e9: data_out = 12'h003;
            11'h01ea: data_out = 12'h202;
            11'h01eb: data_out = 12'h92b;
            11'h01ec: data_out = 12'h220;
            11'h01ed: data_out = 12'h101;
            11'h01ee: data_out = 12'h003;
            11'h01ef: data_out = 12'h202;
            11'h01f0: data_out = 12'h99e;
            11'h01f1: data_out = 12'h221;
            11'h01f2: data_out = 12'h101;
            11'h01f3: data_out = 12'h003;
            11'h01f4: data_out = 12'h202;
            11'h01f5: data_out = 12'h99e;
            11'h01f6: data_out = 12'h230;
            11'h01f7: data_out = 12'h101;
            11'h01f8: data_out = 12'h003;
            11'h01f9: data_out = 12'h203;
            11'h01fa: data_out = 12'h90d;
            11'h01fb: data_out = 12'h231;
            11'h01fc: data_out = 12'h101;
            11'h01fd: data_out = 12'h003;
            11'h01fe: data_out = 12'h203;
            11'h01ff: data_out = 12'h90d;
            11'h0200: data_out = 12'h240;
            11'h0201: data_out = 12'h101;
            11'h0202: data_out = 12'h003;
            11'h0203: data_out = 12'h202;
            11'h0204: data_out = 12'h99a;
            11'h0205: data_out = 12'h241;
            11'h0206: data_out = 12'h101;
            11'h0207: data_out = 12'h003;
            11'h0208: data_out = 12'h202;
            11'h0209: data_out = 12'h99a;
            11'h020a: data_out = 12'h2c4;
            11'h020b: data_out = 12'h101;
            11'h020c: data_out = 12'h003;
            11'h020d: data_out = 12'h202;
            11'h020e: data_out = 12'h99e;
            11'h020f: data_out = 12'h2c5;
            11'h0210: data_out = 12'h101;
            11'h0211: data_out = 12'h003;
            11'h0212: data_out = 12'h203;
            11'h0213: data_out = 12'h90d;
            11'h0214: data_out = 12'h2c6;
            11'h0215: data_out = 12'h101;
            11'h0216: data_out = 12'h003;
            11'h0217: data_out = 12'h202;
            11'h0218: data_out = 12'h923;
            11'h0219: data_out = 12'h270;
            11'h021a: data_out = 12'h101;
            11'h021b: data_out = 12'h003;
            11'h021c: data_out = 12'h201;
            11'h021d: data_out = 12'h9af;
            11'h021e: data_out = 12'h2ec;
            11'h021f: data_out = 12'h101;
            11'h0220: data_out = 12'h003;
            11'h0221: data_out = 12'h203;
            11'h0222: data_out = 12'h969;
            11'h0223: data_out = 12'h201;
            11'h0224: data_out = 12'h100;
            11'h0225: data_out = 12'h205;
            11'h0226: data_out = 12'h4e2;
            11'h0227: data_out = 12'h204;
            11'h0228: data_out = 12'h1c4;
            11'h0229: data_out = 12'h201;
            11'h022a: data_out = 12'h8af;
            11'h022b: data_out = 12'h200;
            11'h022c: data_out = 12'h100;
            11'h022d: data_out = 12'h220;
            11'h022e: data_out = 12'h103;
            11'h022f: data_out = 12'h0c6;
            11'h0230: data_out = 12'h101;
            11'h0231: data_out = 12'h003;
            11'h0232: data_out = 12'h202;
            11'h0233: data_out = 12'h923;
            11'h0234: data_out = 12'h0ca;
            11'h0235: data_out = 12'h101;
            11'h0236: data_out = 12'h003;
            11'h0237: data_out = 12'h202;
            11'h0238: data_out = 12'h923;
            11'h0239: data_out = 12'h0c6;
            11'h023a: data_out = 12'h197;
            11'h023b: data_out = 12'h0ca;
            11'h023c: data_out = 12'h196;
            11'h023d: data_out = 12'h200;
            11'h023e: data_out = 12'h104;
            11'h023f: data_out = 12'h105;
            11'h0240: data_out = 12'h194;
            11'h0241: data_out = 12'h195;
            11'h0242: data_out = 12'h004;
            11'h0243: data_out = 12'h100;
            11'h0244: data_out = 12'h097;
            11'h0245: data_out = 12'h101;
            11'h0246: data_out = 12'h280;
            11'h0247: data_out = 12'h103;
            11'h0248: data_out = 12'h003;
            11'h0249: data_out = 12'h104;
            11'h024a: data_out = 12'h005;
            11'h024b: data_out = 12'h100;
            11'h024c: data_out = 12'h200;
            11'h024d: data_out = 12'h101;
            11'h024e: data_out = 12'h281;
            11'h024f: data_out = 12'h103;
            11'h0250: data_out = 12'h003;
            11'h0251: data_out = 12'h105;
            11'h0252: data_out = 12'h096;
            11'h0253: data_out = 12'h100;
            11'h0254: data_out = 12'h201;
            11'h0255: data_out = 12'h101;
            11'h0256: data_out = 12'h282;
            11'h0257: data_out = 12'h103;
            11'h0258: data_out = 12'h003;
            11'h0259: data_out = 12'h196;
            11'h025a: data_out = 12'h202;
            11'h025b: data_out = 12'h95e;
            11'h025c: data_out = 12'h202;
            11'h025d: data_out = 12'h842;
            11'h025e: data_out = 12'h0ca;
            11'h025f: data_out = 12'h196;
            11'h0260: data_out = 12'h08c;
            11'h0261: data_out = 12'h186;
            11'h0262: data_out = 12'h08d;
            11'h0263: data_out = 12'h187;
            11'h0264: data_out = 12'h08e;
            11'h0265: data_out = 12'h188;
            11'h0266: data_out = 12'h08f;
            11'h0267: data_out = 12'h189;
            11'h0268: data_out = 12'h086;
            11'h0269: data_out = 12'h100;
            11'h026a: data_out = 12'h004;
            11'h026b: data_out = 12'h101;
            11'h026c: data_out = 12'h282;
            11'h026d: data_out = 12'h103;
            11'h026e: data_out = 12'h003;
            11'h026f: data_out = 12'h186;
            11'h0270: data_out = 12'h087;
            11'h0271: data_out = 12'h100;
            11'h0272: data_out = 12'h005;
            11'h0273: data_out = 12'h101;
            11'h0274: data_out = 12'h283;
            11'h0275: data_out = 12'h103;
            11'h0276: data_out = 12'h003;
            11'h0277: data_out = 12'h187;
            11'h0278: data_out = 12'h200;
            11'h0279: data_out = 12'h101;
            11'h027a: data_out = 12'h088;
            11'h027b: data_out = 12'h100;
            11'h027c: data_out = 12'h003;
            11'h027d: data_out = 12'h188;
            11'h027e: data_out = 12'h089;
            11'h027f: data_out = 12'h100;
            11'h0280: data_out = 12'h003;
            11'h0281: data_out = 12'h189;
            11'h0282: data_out = 12'h202;
            11'h0283: data_out = 12'ha86;
            11'h0284: data_out = 12'h202;
            11'h0285: data_out = 12'h898;
            11'h0286: data_out = 12'h094;
            11'h0287: data_out = 12'h100;
            11'h0288: data_out = 12'h201;
            11'h0289: data_out = 12'h101;
            11'h028a: data_out = 12'h280;
            11'h028b: data_out = 12'h103;
            11'h028c: data_out = 12'h003;
            11'h028d: data_out = 12'h194;
            11'h028e: data_out = 12'h095;
            11'h028f: data_out = 12'h100;
            11'h0290: data_out = 12'h200;
            11'h0291: data_out = 12'h101;
            11'h0292: data_out = 12'h281;
            11'h0293: data_out = 12'h103;
            11'h0294: data_out = 12'h003;
            11'h0295: data_out = 12'h195;
            11'h0296: data_out = 12'h202;
            11'h0297: data_out = 12'h868;
            11'h0298: data_out = 12'h201;
            11'h0299: data_out = 12'h8af;
            11'h029a: data_out = 12'h208;
            11'h029b: data_out = 12'h100;
            11'h029c: data_out = 12'h205;
            11'h029d: data_out = 12'h4d4;
            11'h029e: data_out = 12'h205;
            11'h029f: data_out = 12'h40d;
            11'h02a0: data_out = 12'h2ff;
            11'h02a1: data_out = 12'h180;
            11'h02a2: data_out = 12'h205;
            11'h02a3: data_out = 12'h4f0;
            11'h02a4: data_out = 12'h251;
            11'h02a5: data_out = 12'h180;
            11'h02a6: data_out = 12'h205;
            11'h02a7: data_out = 12'h4f0;
            11'h02a8: data_out = 12'h206;
            11'h02a9: data_out = 12'h454;
            11'h02aa: data_out = 12'h20a;
            11'h02ab: data_out = 12'h104;
            11'h02ac: data_out = 12'h206;
            11'h02ad: data_out = 12'h41e;
            11'h02ae: data_out = 12'h005;
            11'h02af: data_out = 12'h100;
            11'h02b0: data_out = 12'h200;
            11'h02b1: data_out = 12'h101;
            11'h02b2: data_out = 12'h240;
            11'h02b3: data_out = 12'h103;
            11'h02b4: data_out = 12'h003;
            11'h02b5: data_out = 12'h202;
            11'h02b6: data_out = 12'h9b9;
            11'h02b7: data_out = 12'h203;
            11'h02b8: data_out = 12'h801;
            11'h02b9: data_out = 12'h2ff;
            11'h02ba: data_out = 12'h107;
            11'h02bb: data_out = 12'h2ff;
            11'h02bc: data_out = 12'h104;
            11'h02bd: data_out = 12'h2fe;
            11'h02be: data_out = 12'h105;
            11'h02bf: data_out = 12'h206;
            11'h02c0: data_out = 12'h439;
            11'h02c1: data_out = 12'h006;
            11'h02c2: data_out = 12'h100;
            11'h02c3: data_out = 12'h2fe;
            11'h02c4: data_out = 12'h101;
            11'h02c5: data_out = 12'h240;
            11'h02c6: data_out = 12'h103;
            11'h02c7: data_out = 12'h003;
            11'h02c8: data_out = 12'h202;
            11'h02c9: data_out = 12'h9d6;
            11'h02ca: data_out = 12'h007;
            11'h02cb: data_out = 12'h100;
            11'h02cc: data_out = 12'h201;
            11'h02cd: data_out = 12'h101;
            11'h02ce: data_out = 12'h282;
            11'h02cf: data_out = 12'h103;
            11'h02d0: data_out = 12'h003;
            11'h02d1: data_out = 12'h107;
            11'h02d2: data_out = 12'h203;
            11'h02d3: data_out = 12'h901;
            11'h02d4: data_out = 12'h202;
            11'h02d5: data_out = 12'h8bb;
            11'h02d6: data_out = 12'h2ff;
            11'h02d7: data_out = 12'h104;
            11'h02d8: data_out = 12'h201;
            11'h02d9: data_out = 12'h105;
            11'h02da: data_out = 12'h2ff;
            11'h02db: data_out = 12'h180;
            11'h02dc: data_out = 12'h205;
            11'h02dd: data_out = 12'h4f0;
            11'h02de: data_out = 12'h080;
            11'h02df: data_out = 12'h1c1;
            11'h02e0: data_out = 12'h206;
            11'h02e1: data_out = 12'h48d;
            11'h02e2: data_out = 12'h202;
            11'h02e3: data_out = 12'hada;
            11'h02e4: data_out = 12'h204;
            11'h02e5: data_out = 12'h4fd;
            11'h02e6: data_out = 12'h082;
            11'h02e7: data_out = 12'h100;
            11'h02e8: data_out = 12'h208;
            11'h02e9: data_out = 12'h101;
            11'h02ea: data_out = 12'h200;
            11'h02eb: data_out = 12'h103;
            11'h02ec: data_out = 12'h003;
            11'h02ed: data_out = 12'h202;
            11'h02ee: data_out = 12'h9f1;
            11'h02ef: data_out = 12'h202;
            11'h02f0: data_out = 12'h8f3;
            11'h02f1: data_out = 12'h205;
            11'h02f2: data_out = 12'h4c0;
            11'h02f3: data_out = 12'h0c6;
            11'h02f4: data_out = 12'h100;
            11'h02f5: data_out = 12'h201;
            11'h02f6: data_out = 12'h101;
            11'h02f7: data_out = 12'h282;
            11'h02f8: data_out = 12'h103;
            11'h02f9: data_out = 12'h003;
            11'h02fa: data_out = 12'h1c6;
            11'h02fb: data_out = 12'h203;
            11'h02fc: data_out = 12'h907;
            11'h02fd: data_out = 12'h205;
            11'h02fe: data_out = 12'h4a7;
            11'h02ff: data_out = 12'h202;
            11'h0300: data_out = 12'h8a0;
            11'h0301: data_out = 12'h240;
            11'h0302: data_out = 12'h1c4;
            11'h0303: data_out = 12'h201;
            11'h0304: data_out = 12'h100;
            11'h0305: data_out = 12'h205;
            11'h0306: data_out = 12'h405;
            11'h0307: data_out = 12'h0f7;
            11'h0308: data_out = 12'h100;
            11'h0309: data_out = 12'h205;
            11'h030a: data_out = 12'h4db;
            11'h030b: data_out = 12'h201;
            11'h030c: data_out = 12'h8af;
            11'h030d: data_out = 12'h205;
            11'h030e: data_out = 12'h40d;
            11'h030f: data_out = 12'h205;
            11'h0310: data_out = 12'h4c0;
            11'h0311: data_out = 12'h2ff;
            11'h0312: data_out = 12'h180;
            11'h0313: data_out = 12'h205;
            11'h0314: data_out = 12'h4f0;
            11'h0315: data_out = 12'h258;
            11'h0316: data_out = 12'h180;
            11'h0317: data_out = 12'h205;
            11'h0318: data_out = 12'h4f0;
            11'h0319: data_out = 12'h206;
            11'h031a: data_out = 12'h454;
            11'h031b: data_out = 12'h20a;
            11'h031c: data_out = 12'h104;
            11'h031d: data_out = 12'h206;
            11'h031e: data_out = 12'h41e;
            11'h031f: data_out = 12'h005;
            11'h0320: data_out = 12'h100;
            11'h0321: data_out = 12'h200;
            11'h0322: data_out = 12'h101;
            11'h0323: data_out = 12'h240;
            11'h0324: data_out = 12'h103;
            11'h0325: data_out = 12'h003;
            11'h0326: data_out = 12'h203;
            11'h0327: data_out = 12'h92a;
            11'h0328: data_out = 12'h203;
            11'h0329: data_out = 12'h861;
            11'h032a: data_out = 12'h2ff;
            11'h032b: data_out = 12'h104;
            11'h032c: data_out = 12'h201;
            11'h032d: data_out = 12'h105;
            11'h032e: data_out = 12'h2ff;
            11'h032f: data_out = 12'h180;
            11'h0330: data_out = 12'h205;
            11'h0331: data_out = 12'h4f0;
            11'h0332: data_out = 12'h2fe;
            11'h0333: data_out = 12'h180;
            11'h0334: data_out = 12'h205;
            11'h0335: data_out = 12'h4f0;
            11'h0336: data_out = 12'h0c1;
            11'h0337: data_out = 12'h180;
            11'h0338: data_out = 12'h205;
            11'h0339: data_out = 12'h4f0;
            11'h033a: data_out = 12'h206;
            11'h033b: data_out = 12'h48d;
            11'h033c: data_out = 12'h203;
            11'h033d: data_out = 12'ha36;
            11'h033e: data_out = 12'h206;
            11'h033f: data_out = 12'h400;
            11'h0340: data_out = 12'h080;
            11'h0341: data_out = 12'h100;
            11'h0342: data_out = 12'h21f;
            11'h0343: data_out = 12'h101;
            11'h0344: data_out = 12'h200;
            11'h0345: data_out = 12'h103;
            11'h0346: data_out = 12'h003;
            11'h0347: data_out = 12'h100;
            11'h0348: data_out = 12'h205;
            11'h0349: data_out = 12'h101;
            11'h034a: data_out = 12'h240;
            11'h034b: data_out = 12'h103;
            11'h034c: data_out = 12'h003;
            11'h034d: data_out = 12'h203;
            11'h034e: data_out = 12'h951;
            11'h034f: data_out = 12'h203;
            11'h0350: data_out = 12'h861;
            11'h0351: data_out = 12'h204;
            11'h0352: data_out = 12'h4fd;
            11'h0353: data_out = 12'h0c6;
            11'h0354: data_out = 12'h100;
            11'h0355: data_out = 12'h201;
            11'h0356: data_out = 12'h101;
            11'h0357: data_out = 12'h282;
            11'h0358: data_out = 12'h103;
            11'h0359: data_out = 12'h003;
            11'h035a: data_out = 12'h1c6;
            11'h035b: data_out = 12'h203;
            11'h035c: data_out = 12'h967;
            11'h035d: data_out = 12'h205;
            11'h035e: data_out = 12'h4a7;
            11'h035f: data_out = 12'h203;
            11'h0360: data_out = 12'h80f;
            11'h0361: data_out = 12'h240;
            11'h0362: data_out = 12'h1c4;
            11'h0363: data_out = 12'h201;
            11'h0364: data_out = 12'h100;
            11'h0365: data_out = 12'h205;
            11'h0366: data_out = 12'h405;
            11'h0367: data_out = 12'h201;
            11'h0368: data_out = 12'h8af;
            11'h0369: data_out = 12'h240;
            11'h036a: data_out = 12'h1c1;
            11'h036b: data_out = 12'h200;
            11'h036c: data_out = 12'h1c1;
            11'h036d: data_out = 12'h090;
            11'h036e: data_out = 12'h1c1;
            11'h036f: data_out = 12'h091;
            11'h0370: data_out = 12'h1c1;
            11'h0371: data_out = 12'h200;
            11'h0372: data_out = 12'h1c1;
            11'h0373: data_out = 12'h200;
            11'h0374: data_out = 12'h1c1;
            11'h0375: data_out = 12'h092;
            11'h0376: data_out = 12'h1c1;
            11'h0377: data_out = 12'h200;
            11'h0378: data_out = 12'h1c1;
            11'h0379: data_out = 12'h200;
            11'h037a: data_out = 12'h1c1;
            11'h037b: data_out = 12'h200;
            11'h037c: data_out = 12'h1c1;
            11'h037d: data_out = 12'h200;
            11'h037e: data_out = 12'h1c1;
            11'h037f: data_out = 12'h200;
            11'h0380: data_out = 12'h1c1;
            11'h0381: data_out = 12'h093;
            11'h0382: data_out = 12'h1c1;
            11'h0383: data_out = 12'h200;
            11'h0384: data_out = 12'h1c1;
            11'h0385: data_out = 12'h200;
            11'h0386: data_out = 12'h1c1;
            11'h0387: data_out = 12'h200;
            11'h0388: data_out = 12'h1c1;
            11'h0389: data_out = 12'h200;
            11'h038a: data_out = 12'h1c1;
            11'h038b: data_out = 12'h200;
            11'h038c: data_out = 12'h1c1;
            11'h038d: data_out = 12'h200;
            11'h038e: data_out = 12'h1c1;
            11'h038f: data_out = 12'h200;
            11'h0390: data_out = 12'h1c1;
            11'h0391: data_out = 12'h246;
            11'h0392: data_out = 12'h1c1;
            11'h0393: data_out = 12'h24b;
            11'h0394: data_out = 12'h1c1;
            11'h0395: data_out = 12'h24d;
            11'h0396: data_out = 12'h1c1;
            11'h0397: data_out = 12'h24d;
            11'h0398: data_out = 12'h1c1;
            11'h0399: data_out = 12'h249;
            11'h039a: data_out = 12'h1c1;
            11'h039b: data_out = 12'h243;
            11'h039c: data_out = 12'h1c1;
            11'h039d: data_out = 12'h245;
            11'h039e: data_out = 12'h1c1;
            11'h039f: data_out = 12'h244;
            11'h03a0: data_out = 12'h1c1;
            11'h03a1: data_out = 12'h230;
            11'h03a2: data_out = 12'h1c1;
            11'h03a3: data_out = 12'h230;
            11'h03a4: data_out = 12'h1c1;
            11'h03a5: data_out = 12'h230;
            11'h03a6: data_out = 12'h1c1;
            11'h03a7: data_out = 12'h230;
            11'h03a8: data_out = 12'h1c1;
            11'h03a9: data_out = 12'h220;
            11'h03aa: data_out = 12'h1c1;
            11'h03ab: data_out = 12'h230;
            11'h03ac: data_out = 12'h1c1;
            11'h03ad: data_out = 12'h220;
            11'h03ae: data_out = 12'h1c1;
            11'h03af: data_out = 12'h220;
            11'h03b0: data_out = 12'h1c1;
            11'h03b1: data_out = 12'h220;
            11'h03b2: data_out = 12'h1c1;
            11'h03b3: data_out = 12'h220;
            11'h03b4: data_out = 12'h1c1;
            11'h03b5: data_out = 12'h220;
            11'h03b6: data_out = 12'h1c1;
            11'h03b7: data_out = 12'h220;
            11'h03b8: data_out = 12'h1c1;
            11'h03b9: data_out = 12'h200;
            11'h03ba: data_out = 12'h1c1;
            11'h03bb: data_out = 12'h200;
            11'h03bc: data_out = 12'h1c1;
            11'h03bd: data_out = 12'h200;
            11'h03be: data_out = 12'h1c1;
            11'h03bf: data_out = 12'h200;
            11'h03c0: data_out = 12'h1c1;
            11'h03c1: data_out = 12'h200;
            11'h03c2: data_out = 12'h1c1;
            11'h03c3: data_out = 12'h200;
            11'h03c4: data_out = 12'h1c1;
            11'h03c5: data_out = 12'h230;
            11'h03c6: data_out = 12'h1c1;
            11'h03c7: data_out = 12'h230;
            11'h03c8: data_out = 12'h1c1;
            11'h03c9: data_out = 12'h230;
            11'h03ca: data_out = 12'h1c1;
            11'h03cb: data_out = 12'h230;
            11'h03cc: data_out = 12'h1c1;
            11'h03cd: data_out = 12'h230;
            11'h03ce: data_out = 12'h1c1;
            11'h03cf: data_out = 12'h230;
            11'h03d0: data_out = 12'h1c1;
            11'h03d1: data_out = 12'h230;
            11'h03d2: data_out = 12'h1c1;
            11'h03d3: data_out = 12'h230;
            11'h03d4: data_out = 12'h1c1;
            11'h03d5: data_out = 12'h246;
            11'h03d6: data_out = 12'h1c1;
            11'h03d7: data_out = 12'h24b;
            11'h03d8: data_out = 12'h1c1;
            11'h03d9: data_out = 12'h24d;
            11'h03da: data_out = 12'h1c1;
            11'h03db: data_out = 12'h24d;
            11'h03dc: data_out = 12'h1c1;
            11'h03dd: data_out = 12'h249;
            11'h03de: data_out = 12'h1c1;
            11'h03df: data_out = 12'h243;
            11'h03e0: data_out = 12'h1c1;
            11'h03e1: data_out = 12'h245;
            11'h03e2: data_out = 12'h1c1;
            11'h03e3: data_out = 12'h244;
            11'h03e4: data_out = 12'h1c1;
            11'h03e5: data_out = 12'h230;
            11'h03e6: data_out = 12'h1c1;
            11'h03e7: data_out = 12'h230;
            11'h03e8: data_out = 12'h1c1;
            11'h03e9: data_out = 12'h230;
            11'h03ea: data_out = 12'h1c1;
            11'h03eb: data_out = 12'h230;
            11'h03ec: data_out = 12'h1c1;
            11'h03ed: data_out = 12'h220;
            11'h03ee: data_out = 12'h1c1;
            11'h03ef: data_out = 12'h230;
            11'h03f0: data_out = 12'h1c1;
            11'h03f1: data_out = 12'h220;
            11'h03f2: data_out = 12'h1c1;
            11'h03f3: data_out = 12'h220;
            11'h03f4: data_out = 12'h1c1;
            11'h03f5: data_out = 12'h220;
            11'h03f6: data_out = 12'h1c1;
            11'h03f7: data_out = 12'h220;
            11'h03f8: data_out = 12'h1c1;
            11'h03f9: data_out = 12'h220;
            11'h03fa: data_out = 12'h1c1;
            11'h03fb: data_out = 12'h220;
            11'h03fc: data_out = 12'h1c1;
            11'h03fd: data_out = 12'h220;
            11'h03fe: data_out = 12'h1c1;
            11'h03ff: data_out = 12'h220;
            11'h0400: data_out = 12'h1c1;
            11'h0401: data_out = 12'h220;
            11'h0402: data_out = 12'h1c1;
            11'h0403: data_out = 12'h220;
            11'h0404: data_out = 12'h1c1;
            11'h0405: data_out = 12'h220;
            11'h0406: data_out = 12'h1c1;
            11'h0407: data_out = 12'h220;
            11'h0408: data_out = 12'h1c1;
            11'h0409: data_out = 12'h220;
            11'h040a: data_out = 12'h1c1;
            11'h040b: data_out = 12'h220;
            11'h040c: data_out = 12'h1c1;
            11'h040d: data_out = 12'h220;
            11'h040e: data_out = 12'h1c1;
            11'h040f: data_out = 12'h220;
            11'h0410: data_out = 12'h1c1;
            11'h0411: data_out = 12'h220;
            11'h0412: data_out = 12'h1c1;
            11'h0413: data_out = 12'h220;
            11'h0414: data_out = 12'h1c1;
            11'h0415: data_out = 12'h220;
            11'h0416: data_out = 12'h1c1;
            11'h0417: data_out = 12'h220;
            11'h0418: data_out = 12'h1c1;
            11'h0419: data_out = 12'h220;
            11'h041a: data_out = 12'h1c1;
            11'h041b: data_out = 12'h220;
            11'h041c: data_out = 12'h1c1;
            11'h041d: data_out = 12'h220;
            11'h041e: data_out = 12'h1c1;
            11'h041f: data_out = 12'h220;
            11'h0420: data_out = 12'h1c1;
            11'h0421: data_out = 12'h220;
            11'h0422: data_out = 12'h1c1;
            11'h0423: data_out = 12'h220;
            11'h0424: data_out = 12'h1c1;
            11'h0425: data_out = 12'h201;
            11'h0426: data_out = 12'h1c1;
            11'h0427: data_out = 12'h280;
            11'h0428: data_out = 12'h1c1;
            11'h0429: data_out = 12'h200;
            11'h042a: data_out = 12'h1c1;
            11'h042b: data_out = 12'h200;
            11'h042c: data_out = 12'h1c1;
            11'h042d: data_out = 12'h200;
            11'h042e: data_out = 12'h1c1;
            11'h042f: data_out = 12'h202;
            11'h0430: data_out = 12'h1c1;
            11'h0431: data_out = 12'h201;
            11'h0432: data_out = 12'h1c1;
            11'h0433: data_out = 12'h240;
            11'h0434: data_out = 12'h1c1;
            11'h0435: data_out = 12'h200;
            11'h0436: data_out = 12'h1c1;
            11'h0437: data_out = 12'h202;
            11'h0438: data_out = 12'h1c1;
            11'h0439: data_out = 12'h200;
            11'h043a: data_out = 12'h1c1;
            11'h043b: data_out = 12'h202;
            11'h043c: data_out = 12'h1c1;
            11'h043d: data_out = 12'h207;
            11'h043e: data_out = 12'h1c1;
            11'h043f: data_out = 12'h200;
            11'h0440: data_out = 12'h1c1;
            11'h0441: data_out = 12'h094;
            11'h0442: data_out = 12'h1c1;
            11'h0443: data_out = 12'h095;
            11'h0444: data_out = 12'h1c1;
            11'h0445: data_out = 12'h096;
            11'h0446: data_out = 12'h1c1;
            11'h0447: data_out = 12'h200;
            11'h0448: data_out = 12'h1c1;
            11'h0449: data_out = 12'h097;
            11'h044a: data_out = 12'h1c1;
            11'h044b: data_out = 12'h200;
            11'h044c: data_out = 12'h1c1;
            11'h044d: data_out = 12'h08c;
            11'h044e: data_out = 12'h1c1;
            11'h044f: data_out = 12'h08d;
            11'h0450: data_out = 12'h1c1;
            11'h0451: data_out = 12'h08e;
            11'h0452: data_out = 12'h1c1;
            11'h0453: data_out = 12'h08f;
            11'h0454: data_out = 12'h1c1;
            11'h0455: data_out = 12'h200;
            11'h0456: data_out = 12'h1c1;
            11'h0457: data_out = 12'h200;
            11'h0458: data_out = 12'h1c1;
            11'h0459: data_out = 12'h08c;
            11'h045a: data_out = 12'h1c1;
            11'h045b: data_out = 12'h08d;
            11'h045c: data_out = 12'h1c1;
            11'h045d: data_out = 12'h08e;
            11'h045e: data_out = 12'h1c1;
            11'h045f: data_out = 12'h08f;
            11'h0460: data_out = 12'h1c1;
            11'h0461: data_out = 12'h200;
            11'h0462: data_out = 12'h1c1;
            11'h0463: data_out = 12'h200;
            11'h0464: data_out = 12'h1c1;
            11'h0465: data_out = 12'h200;
            11'h0466: data_out = 12'h1c1;
            11'h0467: data_out = 12'h200;
            11'h0468: data_out = 12'h1c1;
            11'h0469: data_out = 12'h200;
            11'h046a: data_out = 12'h1c1;
            11'h046b: data_out = 12'h200;
            11'h046c: data_out = 12'h1c1;
            11'h046d: data_out = 12'h278;
            11'h046e: data_out = 12'h1c1;
            11'h046f: data_out = 12'h200;
            11'h0470: data_out = 12'h1c1;
            11'h0471: data_out = 12'h278;
            11'h0472: data_out = 12'h1c1;
            11'h0473: data_out = 12'h200;
            11'h0474: data_out = 12'h1c1;
            11'h0475: data_out = 12'h278;
            11'h0476: data_out = 12'h1c1;
            11'h0477: data_out = 12'h200;
            11'h0478: data_out = 12'h1c1;
            11'h0479: data_out = 12'h278;
            11'h047a: data_out = 12'h1c1;
            11'h047b: data_out = 12'h200;
            11'h047c: data_out = 12'h1c1;
            11'h047d: data_out = 12'h200;
            11'h047e: data_out = 12'h1c1;
            11'h047f: data_out = 12'h200;
            11'h0480: data_out = 12'h1c1;
            11'h0481: data_out = 12'h200;
            11'h0482: data_out = 12'h1c1;
            11'h0483: data_out = 12'h200;
            11'h0484: data_out = 12'h1c1;
            11'h0485: data_out = 12'h200;
            11'h0486: data_out = 12'h1c1;
            11'h0487: data_out = 12'h200;
            11'h0488: data_out = 12'h1c1;
            11'h0489: data_out = 12'h200;
            11'h048a: data_out = 12'h1c1;
            11'h048b: data_out = 12'h200;
            11'h048c: data_out = 12'h1c1;
            11'h048d: data_out = 12'h200;
            11'h048e: data_out = 12'h1c1;
            11'h048f: data_out = 12'h200;
            11'h0490: data_out = 12'h1c1;
            11'h0491: data_out = 12'h200;
            11'h0492: data_out = 12'h1c1;
            11'h0493: data_out = 12'h200;
            11'h0494: data_out = 12'h1c1;
            11'h0495: data_out = 12'h200;
            11'h0496: data_out = 12'h1c1;
            11'h0497: data_out = 12'h200;
            11'h0498: data_out = 12'h1c1;
            11'h0499: data_out = 12'h200;
            11'h049a: data_out = 12'h1c1;
            11'h049b: data_out = 12'h200;
            11'h049c: data_out = 12'h1c1;
            11'h049d: data_out = 12'h200;
            11'h049e: data_out = 12'h1c1;
            11'h049f: data_out = 12'h200;
            11'h04a0: data_out = 12'h1c1;
            11'h04a1: data_out = 12'h200;
            11'h04a2: data_out = 12'h1c1;
            11'h04a3: data_out = 12'h200;
            11'h04a4: data_out = 12'h1c1;
            11'h04a5: data_out = 12'h200;
            11'h04a6: data_out = 12'h1c1;
            11'h04a7: data_out = 12'h200;
            11'h04a8: data_out = 12'h1c1;
            11'h04a9: data_out = 12'h27e;
            11'h04aa: data_out = 12'h1c1;
            11'h04ab: data_out = 12'h200;
            11'h04ac: data_out = 12'h1c1;
            11'h04ad: data_out = 12'h200;
            11'h04ae: data_out = 12'h1c1;
            11'h04af: data_out = 12'h200;
            11'h04b0: data_out = 12'h1c1;
            11'h04b1: data_out = 12'h200;
            11'h04b2: data_out = 12'h1c1;
            11'h04b3: data_out = 12'h200;
            11'h04b4: data_out = 12'h1c1;
            11'h04b5: data_out = 12'h200;
            11'h04b6: data_out = 12'h1c1;
            11'h04b7: data_out = 12'h200;
            11'h04b8: data_out = 12'h1c1;
            11'h04b9: data_out = 12'h200;
            11'h04ba: data_out = 12'h1c1;
            11'h04bb: data_out = 12'h200;
            11'h04bc: data_out = 12'h1c1;
            11'h04bd: data_out = 12'h200;
            11'h04be: data_out = 12'h1c1;
            11'h04bf: data_out = 12'h200;
            11'h04c0: data_out = 12'h1c1;
            11'h04c1: data_out = 12'h200;
            11'h04c2: data_out = 12'h1c1;
            11'h04c3: data_out = 12'h200;
            11'h04c4: data_out = 12'h1c1;
            11'h04c5: data_out = 12'h200;
            11'h04c6: data_out = 12'h1c1;
            11'h04c7: data_out = 12'h200;
            11'h04c8: data_out = 12'h1c1;
            11'h04c9: data_out = 12'h200;
            11'h04ca: data_out = 12'h1c1;
            11'h04cb: data_out = 12'h200;
            11'h04cc: data_out = 12'h1c1;
            11'h04cd: data_out = 12'h200;
            11'h04ce: data_out = 12'h1c1;
            11'h04cf: data_out = 12'h200;
            11'h04d0: data_out = 12'h1c1;
            11'h04d1: data_out = 12'h200;
            11'h04d2: data_out = 12'h1c1;
            11'h04d3: data_out = 12'h200;
            11'h04d4: data_out = 12'h1c1;
            11'h04d5: data_out = 12'h200;
            11'h04d6: data_out = 12'h1c1;
            11'h04d7: data_out = 12'h200;
            11'h04d8: data_out = 12'h1c1;
            11'h04d9: data_out = 12'h200;
            11'h04da: data_out = 12'h1c1;
            11'h04db: data_out = 12'h200;
            11'h04dc: data_out = 12'h1c1;
            11'h04dd: data_out = 12'h20b;
            11'h04de: data_out = 12'h1c1;
            11'h04df: data_out = 12'h263;
            11'h04e0: data_out = 12'h1c1;
            11'h04e1: data_out = 12'h201;
            11'h04e2: data_out = 12'h101;
            11'h04e3: data_out = 12'h282;
            11'h04e4: data_out = 12'h103;
            11'h04e5: data_out = 12'h245;
            11'h04e6: data_out = 12'h100;
            11'h04e7: data_out = 12'h200;
            11'h04e8: data_out = 12'h1c1;
            11'h04e9: data_out = 12'h003;
            11'h04ea: data_out = 12'h100;
            11'h04eb: data_out = 12'h204;
            11'h04ec: data_out = 12'h9ef;
            11'h04ed: data_out = 12'h204;
            11'h04ee: data_out = 12'h8e7;
            11'h04ef: data_out = 12'h2ff;
            11'h04f0: data_out = 12'h100;
            11'h04f1: data_out = 12'h200;
            11'h04f2: data_out = 12'h1c1;
            11'h04f3: data_out = 12'h003;
            11'h04f4: data_out = 12'h100;
            11'h04f5: data_out = 12'h204;
            11'h04f6: data_out = 12'h9f9;
            11'h04f7: data_out = 12'h204;
            11'h04f8: data_out = 12'h8f1;
            11'h04f9: data_out = 12'h205;
            11'h04fa: data_out = 12'h4c0;
            11'h04fb: data_out = 12'h201;
            11'h04fc: data_out = 12'h8af;
            11'h04fd: data_out = 12'h2ff;
            11'h04fe: data_out = 12'h180;
            11'h04ff: data_out = 12'h205;
            11'h0500: data_out = 12'h4f0;
            11'h0501: data_out = 12'h080;
            11'h0502: data_out = 12'h100;
            11'h0503: data_out = 12'h2ff;
            11'h0504: data_out = 12'h101;
            11'h0505: data_out = 12'h240;
            11'h0506: data_out = 12'h103;
            11'h0507: data_out = 12'h003;
            11'h0508: data_out = 12'h205;
            11'h0509: data_out = 12'h90c;
            11'h050a: data_out = 12'h204;
            11'h050b: data_out = 12'h8fd;
            11'h050c: data_out = 12'h500;
            11'h050d: data_out = 12'h0cc;
            11'h050e: data_out = 12'h100;
            11'h050f: data_out = 12'h201;
            11'h0510: data_out = 12'h101;
            11'h0511: data_out = 12'h200;
            11'h0512: data_out = 12'h103;
            11'h0513: data_out = 12'h003;
            11'h0514: data_out = 12'h205;
            11'h0515: data_out = 12'h91f;
            11'h0516: data_out = 12'h0c7;
            11'h0517: data_out = 12'h186;
            11'h0518: data_out = 12'h0c8;
            11'h0519: data_out = 12'h187;
            11'h051a: data_out = 12'h0c9;
            11'h051b: data_out = 12'h188;
            11'h051c: data_out = 12'h0ca;
            11'h051d: data_out = 12'h189;
            11'h051e: data_out = 12'h500;
            11'h051f: data_out = 12'h200;
            11'h0520: data_out = 12'h186;
            11'h0521: data_out = 12'h187;
            11'h0522: data_out = 12'h188;
            11'h0523: data_out = 12'h189;
            11'h0524: data_out = 12'h105;
            11'h0525: data_out = 12'h106;
            11'h0526: data_out = 12'h0ca;
            11'h0527: data_out = 12'h104;
            11'h0528: data_out = 12'h096;
            11'h0529: data_out = 12'h107;
            11'h052a: data_out = 12'h004;
            11'h052b: data_out = 12'h100;
            11'h052c: data_out = 12'h0c8;
            11'h052d: data_out = 12'h101;
            11'h052e: data_out = 12'h280;
            11'h052f: data_out = 12'h103;
            11'h0530: data_out = 12'h003;
            11'h0531: data_out = 12'h104;
            11'h0532: data_out = 12'h005;
            11'h0533: data_out = 12'h100;
            11'h0534: data_out = 12'h0c9;
            11'h0535: data_out = 12'h101;
            11'h0536: data_out = 12'h281;
            11'h0537: data_out = 12'h103;
            11'h0538: data_out = 12'h003;
            11'h0539: data_out = 12'h105;
            11'h053a: data_out = 12'h006;
            11'h053b: data_out = 12'h100;
            11'h053c: data_out = 12'h000;
            11'h053d: data_out = 12'h101;
            11'h053e: data_out = 12'h003;
            11'h053f: data_out = 12'h106;
            11'h0540: data_out = 12'h007;
            11'h0541: data_out = 12'h100;
            11'h0542: data_out = 12'h201;
            11'h0543: data_out = 12'h101;
            11'h0544: data_out = 12'h282;
            11'h0545: data_out = 12'h103;
            11'h0546: data_out = 12'h003;
            11'h0547: data_out = 12'h107;
            11'h0548: data_out = 12'h205;
            11'h0549: data_out = 12'h94c;
            11'h054a: data_out = 12'h205;
            11'h054b: data_out = 12'h82a;
            11'h054c: data_out = 12'h097;
            11'h054d: data_out = 12'h107;
            11'h054e: data_out = 12'h086;
            11'h054f: data_out = 12'h100;
            11'h0550: data_out = 12'h004;
            11'h0551: data_out = 12'h101;
            11'h0552: data_out = 12'h280;
            11'h0553: data_out = 12'h103;
            11'h0554: data_out = 12'h003;
            11'h0555: data_out = 12'h186;
            11'h0556: data_out = 12'h087;
            11'h0557: data_out = 12'h100;
            11'h0558: data_out = 12'h005;
            11'h0559: data_out = 12'h101;
            11'h055a: data_out = 12'h281;
            11'h055b: data_out = 12'h103;
            11'h055c: data_out = 12'h003;
            11'h055d: data_out = 12'h187;
            11'h055e: data_out = 12'h088;
            11'h055f: data_out = 12'h100;
            11'h0560: data_out = 12'h006;
            11'h0561: data_out = 12'h101;
            11'h0562: data_out = 12'h003;
            11'h0563: data_out = 12'h188;
            11'h0564: data_out = 12'h089;
            11'h0565: data_out = 12'h100;
            11'h0566: data_out = 12'h200;
            11'h0567: data_out = 12'h101;
            11'h0568: data_out = 12'h003;
            11'h0569: data_out = 12'h189;
            11'h056a: data_out = 12'h007;
            11'h056b: data_out = 12'h100;
            11'h056c: data_out = 12'h201;
            11'h056d: data_out = 12'h101;
            11'h056e: data_out = 12'h282;
            11'h056f: data_out = 12'h103;
            11'h0570: data_out = 12'h003;
            11'h0571: data_out = 12'h107;
            11'h0572: data_out = 12'h205;
            11'h0573: data_out = 12'h976;
            11'h0574: data_out = 12'h205;
            11'h0575: data_out = 12'h84e;
            11'h0576: data_out = 12'h086;
            11'h0577: data_out = 12'h100;
            11'h0578: data_out = 12'h0c7;
            11'h0579: data_out = 12'h101;
            11'h057a: data_out = 12'h280;
            11'h057b: data_out = 12'h103;
            11'h057c: data_out = 12'h003;
            11'h057d: data_out = 12'h186;
            11'h057e: data_out = 12'h087;
            11'h057f: data_out = 12'h100;
            11'h0580: data_out = 12'h200;
            11'h0581: data_out = 12'h101;
            11'h0582: data_out = 12'h281;
            11'h0583: data_out = 12'h103;
            11'h0584: data_out = 12'h003;
            11'h0585: data_out = 12'h187;
            11'h0586: data_out = 12'h088;
            11'h0587: data_out = 12'h100;
            11'h0588: data_out = 12'h003;
            11'h0589: data_out = 12'h188;
            11'h058a: data_out = 12'h089;
            11'h058b: data_out = 12'h100;
            11'h058c: data_out = 12'h003;
            11'h058d: data_out = 12'h189;
            11'h058e: data_out = 12'h086;
            11'h058f: data_out = 12'h100;
            11'h0590: data_out = 12'h201;
            11'h0591: data_out = 12'h101;
            11'h0592: data_out = 12'h282;
            11'h0593: data_out = 12'h103;
            11'h0594: data_out = 12'h003;
            11'h0595: data_out = 12'h186;
            11'h0596: data_out = 12'h087;
            11'h0597: data_out = 12'h100;
            11'h0598: data_out = 12'h200;
            11'h0599: data_out = 12'h101;
            11'h059a: data_out = 12'h283;
            11'h059b: data_out = 12'h103;
            11'h059c: data_out = 12'h003;
            11'h059d: data_out = 12'h187;
            11'h059e: data_out = 12'h088;
            11'h059f: data_out = 12'h100;
            11'h05a0: data_out = 12'h003;
            11'h05a1: data_out = 12'h188;
            11'h05a2: data_out = 12'h089;
            11'h05a3: data_out = 12'h100;
            11'h05a4: data_out = 12'h003;
            11'h05a5: data_out = 12'h189;
            11'h05a6: data_out = 12'h500;
            11'h05a7: data_out = 12'h086;
            11'h05a8: data_out = 12'h100;
            11'h05a9: data_out = 12'h201;
            11'h05aa: data_out = 12'h101;
            11'h05ab: data_out = 12'h280;
            11'h05ac: data_out = 12'h103;
            11'h05ad: data_out = 12'h003;
            11'h05ae: data_out = 12'h186;
            11'h05af: data_out = 12'h087;
            11'h05b0: data_out = 12'h100;
            11'h05b1: data_out = 12'h200;
            11'h05b2: data_out = 12'h101;
            11'h05b3: data_out = 12'h281;
            11'h05b4: data_out = 12'h103;
            11'h05b5: data_out = 12'h003;
            11'h05b6: data_out = 12'h187;
            11'h05b7: data_out = 12'h088;
            11'h05b8: data_out = 12'h100;
            11'h05b9: data_out = 12'h003;
            11'h05ba: data_out = 12'h188;
            11'h05bb: data_out = 12'h089;
            11'h05bc: data_out = 12'h100;
            11'h05bd: data_out = 12'h003;
            11'h05be: data_out = 12'h189;
            11'h05bf: data_out = 12'h500;
            11'h05c0: data_out = 12'h201;
            11'h05c1: data_out = 12'h1c2;
            11'h05c2: data_out = 12'h27f;
            11'h05c3: data_out = 12'h100;
            11'h05c4: data_out = 12'h205;
            11'h05c5: data_out = 12'h4e9;
            11'h05c6: data_out = 12'h200;
            11'h05c7: data_out = 12'h103;
            11'h05c8: data_out = 12'h208;
            11'h05c9: data_out = 12'h101;
            11'h05ca: data_out = 12'h0c3;
            11'h05cb: data_out = 12'h100;
            11'h05cc: data_out = 12'h003;
            11'h05cd: data_out = 12'h205;
            11'h05ce: data_out = 12'h9d1;
            11'h05cf: data_out = 12'h205;
            11'h05d0: data_out = 12'h8ca;
            11'h05d1: data_out = 12'h280;
            11'h05d2: data_out = 12'h1c3;
            11'h05d3: data_out = 12'h500;
            11'h05d4: data_out = 12'h082;
            11'h05d5: data_out = 12'h101;
            11'h05d6: data_out = 12'h220;
            11'h05d7: data_out = 12'h103;
            11'h05d8: data_out = 12'h003;
            11'h05d9: data_out = 12'h182;
            11'h05da: data_out = 12'h500;
            11'h05db: data_out = 12'h082;
            11'h05dc: data_out = 12'h101;
            11'h05dd: data_out = 12'h200;
            11'h05de: data_out = 12'h103;
            11'h05df: data_out = 12'h003;
            11'h05e0: data_out = 12'h182;
            11'h05e1: data_out = 12'h500;
            11'h05e2: data_out = 12'h0c3;
            11'h05e3: data_out = 12'h101;
            11'h05e4: data_out = 12'h220;
            11'h05e5: data_out = 12'h103;
            11'h05e6: data_out = 12'h003;
            11'h05e7: data_out = 12'h1c3;
            11'h05e8: data_out = 12'h500;
            11'h05e9: data_out = 12'h0c3;
            11'h05ea: data_out = 12'h101;
            11'h05eb: data_out = 12'h200;
            11'h05ec: data_out = 12'h103;
            11'h05ed: data_out = 12'h003;
            11'h05ee: data_out = 12'h1c3;
            11'h05ef: data_out = 12'h500;
            11'h05f0: data_out = 12'h201;
            11'h05f1: data_out = 12'h101;
            11'h05f2: data_out = 12'h081;
            11'h05f3: data_out = 12'h100;
            11'h05f4: data_out = 12'h200;
            11'h05f5: data_out = 12'h103;
            11'h05f6: data_out = 12'h003;
            11'h05f7: data_out = 12'h205;
            11'h05f8: data_out = 12'h9fb;
            11'h05f9: data_out = 12'h205;
            11'h05fa: data_out = 12'h8f0;
            11'h05fb: data_out = 12'h500;
            11'h05fc: data_out = 12'h2ff;
            11'h05fd: data_out = 12'h180;
            11'h05fe: data_out = 12'h205;
            11'h05ff: data_out = 12'h4f0;
            11'h0600: data_out = 12'h2ff;
            11'h0601: data_out = 12'h180;
            11'h0602: data_out = 12'h205;
            11'h0603: data_out = 12'h4f0;
            11'h0604: data_out = 12'h2ff;
            11'h0605: data_out = 12'h180;
            11'h0606: data_out = 12'h205;
            11'h0607: data_out = 12'h4f0;
            11'h0608: data_out = 12'h2ff;
            11'h0609: data_out = 12'h180;
            11'h060a: data_out = 12'h205;
            11'h060b: data_out = 12'h4f0;
            11'h060c: data_out = 12'h500;
            11'h060d: data_out = 12'h200;
            11'h060e: data_out = 12'h180;
            11'h060f: data_out = 12'h205;
            11'h0610: data_out = 12'h4f0;
            11'h0611: data_out = 12'h200;
            11'h0612: data_out = 12'h180;
            11'h0613: data_out = 12'h205;
            11'h0614: data_out = 12'h4f0;
            11'h0615: data_out = 12'h200;
            11'h0616: data_out = 12'h180;
            11'h0617: data_out = 12'h205;
            11'h0618: data_out = 12'h4f0;
            11'h0619: data_out = 12'h200;
            11'h061a: data_out = 12'h180;
            11'h061b: data_out = 12'h205;
            11'h061c: data_out = 12'h4f0;
            11'h061d: data_out = 12'h500;
            11'h061e: data_out = 12'h2ff;
            11'h061f: data_out = 12'h180;
            11'h0620: data_out = 12'h205;
            11'h0621: data_out = 12'h4f0;
            11'h0622: data_out = 12'h080;
            11'h0623: data_out = 12'h105;
            11'h0624: data_out = 12'h100;
            11'h0625: data_out = 12'h280;
            11'h0626: data_out = 12'h101;
            11'h0627: data_out = 12'h200;
            11'h0628: data_out = 12'h103;
            11'h0629: data_out = 12'h003;
            11'h062a: data_out = 12'h206;
            11'h062b: data_out = 12'h938;
            11'h062c: data_out = 12'h004;
            11'h062d: data_out = 12'h100;
            11'h062e: data_out = 12'h201;
            11'h062f: data_out = 12'h101;
            11'h0630: data_out = 12'h282;
            11'h0631: data_out = 12'h103;
            11'h0632: data_out = 12'h003;
            11'h0633: data_out = 12'h104;
            11'h0634: data_out = 12'h206;
            11'h0635: data_out = 12'h938;
            11'h0636: data_out = 12'h206;
            11'h0637: data_out = 12'h81e;
            11'h0638: data_out = 12'h500;
            11'h0639: data_out = 12'h2ff;
            11'h063a: data_out = 12'h180;
            11'h063b: data_out = 12'h205;
            11'h063c: data_out = 12'h4f0;
            11'h063d: data_out = 12'h080;
            11'h063e: data_out = 12'h106;
            11'h063f: data_out = 12'h100;
            11'h0640: data_out = 12'h005;
            11'h0641: data_out = 12'h101;
            11'h0642: data_out = 12'h240;
            11'h0643: data_out = 12'h103;
            11'h0644: data_out = 12'h003;
            11'h0645: data_out = 12'h206;
            11'h0646: data_out = 12'h953;
            11'h0647: data_out = 12'h004;
            11'h0648: data_out = 12'h100;
            11'h0649: data_out = 12'h201;
            11'h064a: data_out = 12'h101;
            11'h064b: data_out = 12'h282;
            11'h064c: data_out = 12'h103;
            11'h064d: data_out = 12'h003;
            11'h064e: data_out = 12'h104;
            11'h064f: data_out = 12'h206;
            11'h0650: data_out = 12'h953;
            11'h0651: data_out = 12'h206;
            11'h0652: data_out = 12'h839;
            11'h0653: data_out = 12'h500;
            11'h0654: data_out = 12'h082;
            11'h0655: data_out = 12'h100;
            11'h0656: data_out = 12'h240;
            11'h0657: data_out = 12'h101;
            11'h0658: data_out = 12'h200;
            11'h0659: data_out = 12'h103;
            11'h065a: data_out = 12'h003;
            11'h065b: data_out = 12'h206;
            11'h065c: data_out = 12'h96e;
            11'h065d: data_out = 12'h089;
            11'h065e: data_out = 12'h180;
            11'h065f: data_out = 12'h205;
            11'h0660: data_out = 12'h4f0;
            11'h0661: data_out = 12'h088;
            11'h0662: data_out = 12'h180;
            11'h0663: data_out = 12'h205;
            11'h0664: data_out = 12'h4f0;
            11'h0665: data_out = 12'h087;
            11'h0666: data_out = 12'h180;
            11'h0667: data_out = 12'h205;
            11'h0668: data_out = 12'h4f0;
            11'h0669: data_out = 12'h086;
            11'h066a: data_out = 12'h180;
            11'h066b: data_out = 12'h205;
            11'h066c: data_out = 12'h4f0;
            11'h066d: data_out = 12'h500;
            11'h066e: data_out = 12'h086;
            11'h066f: data_out = 12'h100;
            11'h0670: data_out = 12'h2a0;
            11'h0671: data_out = 12'h103;
            11'h0672: data_out = 12'h003;
            11'h0673: data_out = 12'h104;
            11'h0674: data_out = 12'h087;
            11'h0675: data_out = 12'h100;
            11'h0676: data_out = 12'h2a1;
            11'h0677: data_out = 12'h103;
            11'h0678: data_out = 12'h003;
            11'h0679: data_out = 12'h105;
            11'h067a: data_out = 12'h088;
            11'h067b: data_out = 12'h100;
            11'h067c: data_out = 12'h003;
            11'h067d: data_out = 12'h180;
            11'h067e: data_out = 12'h205;
            11'h067f: data_out = 12'h4f0;
            11'h0680: data_out = 12'h005;
            11'h0681: data_out = 12'h180;
            11'h0682: data_out = 12'h205;
            11'h0683: data_out = 12'h4f0;
            11'h0684: data_out = 12'h004;
            11'h0685: data_out = 12'h180;
            11'h0686: data_out = 12'h205;
            11'h0687: data_out = 12'h4f0;
            11'h0688: data_out = 12'h200;
            11'h0689: data_out = 12'h180;
            11'h068a: data_out = 12'h205;
            11'h068b: data_out = 12'h4f0;
            11'h068c: data_out = 12'h500;
            11'h068d: data_out = 12'h004;
            11'h068e: data_out = 12'h100;
            11'h068f: data_out = 12'h201;
            11'h0690: data_out = 12'h101;
            11'h0691: data_out = 12'h282;
            11'h0692: data_out = 12'h103;
            11'h0693: data_out = 12'h003;
            11'h0694: data_out = 12'h104;
            11'h0695: data_out = 12'h005;
            11'h0696: data_out = 12'h100;
            11'h0697: data_out = 12'h200;
            11'h0698: data_out = 12'h101;
            11'h0699: data_out = 12'h283;
            11'h069a: data_out = 12'h103;
            11'h069b: data_out = 12'h003;
            11'h069c: data_out = 12'h105;
            11'h069d: data_out = 12'h500;
            default: data_out = 12'hxxx;
        endcase
    end
endmodule
